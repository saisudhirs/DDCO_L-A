module and2(c, a);
input a;
output c;
assign c=! a;
endmodule